///////////////////////////////////////////////////////////////////////////////
// Copyright (c) 2021 Intel Corporation
//
// Permission is hereby granted, free of charge, to any person obtaining a
// copy of this software and associated documentation files (the
//"Software"),
// to deal in the Software without restriction, including without limitation
// the rights to use, copy, modify, merge, publish, distribute, sublicense,
// and/or sell copies of the Software, and to permit persons to whom the
// Software is furnished to do so, subject to the following conditions:
//
// The above copyright notice and this permission notice shall be included
//in
// all copies or substantial portions of the Software.
//
// THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
//OR
// IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
// FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL
//THE
// AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
// LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING
// FROM, OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER
// DEALINGS IN THE SOFTWARE.
/////////////////////////////////////////////////////////////////////////////////

module Sigma0 (
	input hash_size,
	input [63:0] in,
	output [63:0] out
	);

wire [63:0] in_rotr2, in_rotr13, in_rotr22; // Rotated input for SHA-256
wire [63:0] in_rotr28, in_rotr34, in_rotr39; // Rotated input for SHA-384/512

assign in_rotr2  = {32'h0, in[1:0], in[31:2]};
assign in_rotr13 = {32'h0, in[12:0], in[31:13]};
assign in_rotr22 = {32'h0, in[21:0], in[31:22]};

assign in_rotr28 = {in[27:0], in[63:28]}; 
assign in_rotr34 = {in[33:0], in[63:34]}; 
assign in_rotr39 = {in[38:0], in[63:39]}; 

assign out = (hash_size==1'b0) ? (in_rotr2 ^ in_rotr13 ^ in_rotr22) : (in_rotr28 ^ in_rotr34 ^ in_rotr39);

endmodule

