package gen_gpo_controls_pkg;

    localparam GPO_1_RST_SRST_BMC_PLD_R_N_BIT_POS = 0;
    localparam GPO_1_RST_RSMRST_PLD_R_N_BIT_POS = 1;
    localparam GPO_1_FM_SPI_PFR_BMC_BT_MASTER_SEL_BIT_POS = 2;
    localparam GPO_1_FM_SPI_PFR_PCH_MASTER_SEL_BIT_POS = 3;
    localparam GPO_1_RELAY1_BLOCK_DISABLE_BIT_POS = 4;
    localparam GPO_1_RELAY1_FILTER_DISABLE_BIT_POS = 5;
    localparam GPO_1_RELAY2_BLOCK_DISABLE_BIT_POS = 6;
    localparam GPO_1_RELAY2_FILTER_DISABLE_BIT_POS = 7;
    localparam GPO_1_RELAY3_BLOCK_DISABLE_BIT_POS = 8;
    localparam GPO_1_RELAY3_FILTER_DISABLE_BIT_POS = 9;
    localparam GPO_1_PWRGD_DSW_PWROK_R_BIT_POS = 10;
    localparam GPO_1_RST_PFR_EXTRST_N_BIT_POS = 11;
    localparam GPO_1_SPI_MASTER_BMC_PCHN_BIT_POS = 12;
    localparam GPO_1_BMC_SPI_FILTER_DISABLE_BIT_POS = 13;
    localparam GPO_1_PCH_SPI_FILTER_DISABLE_BIT_POS = 14;
    localparam GPO_1_BMC_SPI_CLEAR_IBB_DETECTED_BIT_POS = 15;
    localparam GPO_1_BMC_SPI_ADDR_MODE_SET_3B_BIT_POS = 16;
    localparam GPO_1_TRIGGER_TOP_SWAP_RESET_BIT_POS = 17;
    localparam GPO_1_FM_PFR_SLP_SUS_N_BIT_POS = 18;
    localparam GPO_1_RST_SPI_PFR_BMC_BOOT_N_BIT_POS = 19;
    localparam GPO_1_RST_SPI_PFR_PCH_N_BIT_POS = 20;
    localparam GPO_1_CLEAR_PLTRST_DETECT_FLAG_BIT_POS = 21;

endpackage
