`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//!  \file      SyncWithDefault.v
//!  \author    amr/carlos.l.bernal@intel.com
//!  \date      Oct 2, 2011
//!  \brief     Input Synchronizer module
//////////////////////////////////////////////////////////////////////////////////
//!  \fn         module SyncWithDefault
//!  \brief      
//////////////////////////////////////////////////////////////////////////////////
module SyncWithDefault #(parameter DEFAULT_OUT = 1'b0)
(
    input        iClk,
    input        iRst_n,
    input        iSignal,
    output    oSyncSignal
);
//////////////////////////////////////////////////////////////////////////////////
// Includes
//////////////////////////////////////////////////////////////////////////////////

//////////////////////////////////////////////////////////////////////////////////
// Defines
//////////////////////////////////////////////////////////////////////////////////

//////////////////////////////////////////////////////////////////////////////////
//Internal Signals
//////////////////////////////////////////////////////////////////////////////////
//!
//reg    [1:0]    rvSyncSignal_d;
reg     rSyncSignal_ff1;
reg 	rSyncSignal_ff2;
//////////////////////////////////////////////////////////////////////////////////
//Continous assigment
//////////////////////////////////////////////////////////////////////////////////
assign    oSyncSignal    = rSyncSignal_ff2;
//////////////////////////////////////////////////////////////////////////////////
//Sequential Section
//////////////////////////////////////////////////////////////////////////////////
always @(posedge iClk or negedge iRst_n)
begin
    if( !iRst_n)
    begin
        rSyncSignal_ff1    <= DEFAULT_OUT;
        rSyncSignal_ff2    <= DEFAULT_OUT;
    end
    else
    begin
        rSyncSignal_ff1   <= iSignal;
        rSyncSignal_ff2 <= rSyncSignal_ff1;
    end
end
//////////////////////////////////////////////////////////////////////////////////
//Combinational Section
//////////////////////////////////////////////////////////////////////////////////
//always @*
//begin
  //  rvSyncSignal_d    = {rvSyncSignal_q[0],iSignal};
//end
//////////////////////////////////////////////////////////////////////////////////
//Instances
//////////////////////////////////////////////////////////////////////////////////

endmodule
//////////////////////////////////////////////////////////////////////////////////