// chip_id_ip.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module chip_id_ip (
		input  wire        clkin,      //  clkin.clk
		input  wire        reset,      //  reset.reset
		output wire        data_valid, // output.valid
		output wire [63:0] chip_id     //       .data
	);

	altchip_id #(
		.DEVICE_FAMILY ("MAX 10"),
		.ID_VALUE      (64'b1101111010101101101111101110111111011110101011011011111011101111),
		.ID_VALUE_STR  ("deadbeefdeadbeef")
	) chip_id_ip_inst (
		.clkin      (clkin),      //  clkin.clk
		.reset      (reset),      //  reset.reset
		.data_valid (data_valid), // output.valid
		.chip_id    (chip_id)     //       .data
	);

endmodule
