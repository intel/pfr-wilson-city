`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//!  \file      Toggle.v
//!  \author    amr/carlos.l.bernal@intel.com
//!  \date      Jun 10, 2011
//!  \brief     Toggle
//////////////////////////////////////////////////////////////////////////////////
//!  \fn         module Toggle
//!  \brief      

//////////////////////////////////////////////////////////////////////////////////
module Toggle
(
    input iClk,
    input iRst,
    input iCE,
    output oTSignal
);
//////////////////////////////////////////////////////////////////////////////////
// Includes
//////////////////////////////////////////////////////////////////////////////////

//////////////////////////////////////////////////////////////////////////////////
// Defines
//////////////////////////////////////////////////////////////////////////////////

//////////////////////////////////////////////////////////////////////////////////
// Internal Signals
//////////////////////////////////////////////////////////////////////////////////
//!
reg rT_d;
reg rT_q;
//////////////////////////////////////////////////////////////////////////////////
// Continous assigments
//////////////////////////////////////////////////////////////////////////////////
assign oTSignal = rT_q;
//////////////////////////////////////////////////////////////////////////////////
// Sequential logic
//////////////////////////////////////////////////////////////////////////////////
always @(posedge iClk or posedge iRst)
begin
    if(iRst)
    begin
        rT_q    <=  1'b0;
    end
    else
    begin
        if(iCE)
        begin
            rT_q    <=  rT_d;
        end
        else
        begin
            rT_q    <=  rT_q;
        end
    end
end
//////////////////////////////////////////////////////////////////////////////////
// Combinational logic
//////////////////////////////////////////////////////////////////////////////////
always @*
begin
    rT_d    =   ~rT_q;
end
//////////////////////////////////////////////////////////////////////////////////
// Instances
//////////////////////////////////////////////////////////////////////////////////


//////////////////////////////////////////////////////////////////////////////////
endmodule
