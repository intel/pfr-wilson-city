`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//!  \file      InputsSyncWithDefault.v
//!  \author    amr/carlos.l.bernal@intel.com
//!  \date      Oct 10, 2011
//!  \brief     Input Signal Synchronizer
//////////////////////////////////////////////////////////////////////////////////
//!  \fn         module InputsSyncWithDefault
//!  \brief      
//////////////////////////////////////////////////////////////////////////////////
module InputsSyncWithDefault
	#(parameter SIZE = 1, DEFAULT_OUT=1'b0)
(
    input               iClk,
    input               iRst_n,
    input   [SIZE-1:0]  ivSync,
    output  [SIZE-1:0]  ovSync
);
//////////////////////////////////////////////////////////////////////////////////
// Includes
//////////////////////////////////////////////////////////////////////////////////

//////////////////////////////////////////////////////////////////////////////////
// Defines
//////////////////////////////////////////////////////////////////////////////////

//////////////////////////////////////////////////////////////////////////////////
// Internal Signals
//////////////////////////////////////////////////////////////////////////////////

//////////////////////////////////////////////////////////////////////////////////
// Continous assigments
//////////////////////////////////////////////////////////////////////////////////


//////////////////////////////////////////////////////////////////////////////////
// Sequential logic
//////////////////////////////////////////////////////////////////////////////////

//////////////////////////////////////////////////////////////////////////////////
// Combinational logic
//////////////////////////////////////////////////////////////////////////////////



//////////////////////////////////////////////////////////////////////////////////
// Instances
//////////////////////////////////////////////////////////////////////////////////
genvar i;
generate
    for (i=0; i<SIZE; i=i+1)
    begin: SyncBlock
    SyncWithDefault #(.DEFAULT_OUT(DEFAULT_OUT)) mISync
    (
        .iClk           (iClk), 
        .iRst_n           (iRst_n), 
        .iSignal        (ivSync[i]), 
        .oSyncSignal    (ovSync[i]) 
    );
    
    end
endgenerate
//////////////////////////////////////////////////////////////////////////////////


endmodule
