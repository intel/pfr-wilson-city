`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
/*!
    \brief      <b>IIC Registers Module</b>\n
    \details    \n
    \file       NeonCityEventsBRAMRegs.v
    \date       Aug 25, 2012
    \brief      $RCSfile: NeonCityEventsBRAMRegs.v.rca $
                $Date: $
                $Author:  $
                $Revision:  $
                $Aliases: $
                $Log: NeonCityEventsBRAMRegs.v.rca $
                
    \copyright Intel Proprietary -- Copyright 2015 Intel -- All rights reserved
    
*/
//////////////////////////////////////////////////////////////////////////////////
module EventsBRAMRegs
(   
    //! Module's clock input
    input           iClk,
    //! Reset input
    input           iRst,
    //! Enable input
    input           iEnable,
    //!
    output          oAccessDone,
    //! App Access
    input   [9:0]   ivAddress,
    input           iAppWE,
    input   [31:0]  ivAppData,
    input           iAppDataRst,    
    //! SMBus regs access
    input   [11:0]   ivRegID,
    output  [7:0]	 ovRegData
);
//////////////////////////////////////////////////////////////////////////////////
// Includes
//////////////////////////////////////////////////////////////////////////////////

//////////////////////////////////////////////////////////////////////////////////
// Defines
//////////////////////////////////////////////////////////////////////////////////

//////////////////////////////////////////////////////////////////////////////////
// Internal Signals
//////////////////////////////////////////////////////////////////////////////////
//!
wire        wDone;
//!
wire    [7:0]   wvRegOutData;
//////////////////////////////////////////////////////////////////////////////////
// Continous assigments
//////////////////////////////////////////////////////////////////////////////////
assign  oAccessDone =   wDone;
assign  ovRegData   =   wvRegOutData;
//////////////////////////////////////////////////////////////////////////////////
// Sequential logic
//////////////////////////////////////////////////////////////////////////////////

//////////////////////////////////////////////////////////////////////////////////
// Combinational logic
//////////////////////////////////////////////////////////////////////////////////

//////////////////////////////////////////////////////////////////////////////////
// Instances
//////////////////////////////////////////////////////////////////////////////////
Mem1Kx32_4Kx8 mEventBRAM
(
    .iClk           ( iClk ),
    .ivAddressA     ( ivAddress ),  //10 bits
    .ivAddressB     ( ivRegID ),    //11 bits
    .iWE            ( iAppWE ),
    .ivData         ( ivAppData ),  //32 bits
    .ovData         ( wvRegOutData ) //8 bits
);
//
//
//
uDelay #
(
    .TOTAL_BITS(4)
) mAccessDoneDelay
(
    .iClk           ( iClk ),
    .iRst           ( iRst ),
    .iCE            ( 1'b1),
    .iSignal        ( iEnable ),
    .oDelayedIn     ( wDone )
);
/////////////////////////////////////////////////////////////////////////////////


endmodule
